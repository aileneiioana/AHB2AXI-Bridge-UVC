//------------------------------------
// File name   : test_lib.sv
// Author      : EASYIC ENG
// Created     : xx.yy.zzzz
// Description :
//------------------------------------

`include "test_base.sv"
`include "test_example_1.sv"
