//------------------------------------
// File name   : axi_types.sv
// Author      : EASYIC ENG
// Created     : xx.yy.zzzz
// Description :
//------------------------------------

`ifndef AXI_TYPES_SV
`define AXI_TYPES_SV

typedef enum bit {AXI_MASTER, AXI_SLAVE } axi_agent_kind_t;


`endif
