//------------------------------------
// File name   : test_lib.sv
// Author      : EASYIC ENG
// Created     : xx.yy.zzzz
// Description :
//-----------------------------------


`include "axi_agent_config.sv"
`include "test_base.sv"
`include "test_example_1.sv"
`include "test_example_2.sv"
`include "test_example_3.sv"
`include "test_example_4.sv"
`include "test_example_5.sv"
`include "test_example_6.sv"
`include "test_example_7.sv"
`include "test_example_8.sv"
`include "test_example_9.sv"
`include "test_example_10.sv"
`include "test_example_11.sv"
`include "test_example_12.sv"